module biss_tb ();


reg     clk ;
reg     rx  ;
reg     rst ;
reg     verify_rx;

wire    syn_biss_clk ;

//对 biss 实例化
biss biss_inst
(
    .clk    (clk )  ,
    .rx     (rx)    ,
    .rst    (rst)   ,
    .verify_rx  (verify_rx), // 此信号在程序中没体现打算作为该程序总控FPGA 同意接收数据
    .syn_biss_clk (syn_biss_clk )   // 输出给编码器的时钟
);

// 初始化 赋值
initial 
begin
    clk = 0 ;
    rx  = 0 ;
    rst = 0 ;
    verify_rx = 0;   

    #100
    rst = 1;
    verify_rx = 1;

    #1300
    rx = 1 ; //编码器准备好
    #3294
    rx  = 0 ;// 编码器做出应答，低电平输出
    #6578
    rx = 1; // start 位

    #1000
    rx  = 0 ; //0 位
    #1000
    rx  = 1 ; //1 位
    #1000
    rx  = 0 ; //2 位
    #1000
    rx  = 1 ; //3 位
    #1000
    rx  = 0 ; //4 位
    #1000
    rx  = 1 ; //5 位
    #1000
    rx  = 1 ; //6 位
    #1000
    rx  = 0 ; //7 位
    #1000
    rx  = 1 ; //8 位
    #1000
    rx  = 0 ; //9 位
    #1000
    rx  = 1 ; //10 位
    #1000
    rx  = 1 ; //11 位
    #1000
    rx  = 0 ; //12 位
    #1000
    rx  = 1 ; //13 位
    #1000
    rx  = 1 ; //14 位
    #1000
    rx  = 0 ; //15 位
    #1000
    rx  = 1 ; //16 位
    #1000
    rx  = 0 ; //17 位
    #1000
    rx  = 1 ; //18 位
    #1000
    rx  = 1 ; //19 位
    #1000
    rx  = 0 ; //20 位
    #1000
    rx  = 0 ; //21 位
    #1000
    rx  = 1 ; //22 位
    #1000
    rx  = 1 ; //23 位
    #1000
    rx  = 0 ; //24 位
    #1000
    rx  = 1 ; //25 位
    #1000
    rx  = 1 ; //26 位
    #1000
    rx  = 1 ; //27 位 error
    #1000
    rx  = 0 ; //28  warn 位
    #1000
    rx  = 0 ; //29 crc 1 位
    #1000
    rx  = 0 ; //30 crc 2 位
    #1000
    rx  = 0 ; //31 crc 3 位
    #1000
    rx  = 0 ; //32 crc 4 位
    #1000
    rx  = 0 ; //33 crc 5 位
    #1000
    rx  = 0 ; //34 crc 6 位
    #1000
    rx  = 0 ; // 编码器持续输出 低电平
    
   //第二组数据
		#1300
		rx = 1;//编码器输出准备好
		#5764
		rx = 0;//编码器做出应答，低电平输出
		#6893
		rx = 1;//start位
		#1000
		rx = 0;//0位
		#1000
		rx = 1;//1
		#1000
		rx = 0;//2位		
		#1000
		rx = 1;//3位	
		#1000
		rx = 0;//4位	
		#1000
		rx = 1;//5位
		#1000
		rx = 1;//6位
		#1000
		rx = 0;//7位
		#1000
		rx = 1;//8位
		#1000
		rx = 0;//9位
		#1000
		rx = 1;//10位
		#1000
		rx = 1;//11位
		#1000
		rx = 0;//12位
		#1000
		rx = 1;//13位
		#1000
		rx = 1;//14位
		#1000
		rx = 0;//15位
		#1000
		rx = 1;//16位
		#1000
		rx = 0;//17位
		#1000
		rx = 1;//18位
		#1000
		rx = 1;//19位
		#1000
		rx = 0;//20位
		#1000
		rx = 0;//21位
		#1000
		rx = 1;//22位
		#1000
		rx = 1;//23位
		#1000
		rx = 0;//24位
		#1000
		rx = 1;//25位
		#1000
		rx = 1;//26位
		#1000
		rx = 1;//Error，27
		#1000
		rx = 0;//warn位，28
		#1000
		rx = 1;//crc1位，29
		#1000
		rx = 0;//crc2位，30
		#1000
		rx = 1;//crc3位，31
		#1000
		rx = 0;//crc4位，32
		#1000
		rx = 1;//crc5位，33
		#1000
		rx = 1;//crc6位，34
		#1000
		rx = 0;//编码器输出低电平		    


end

// 产生50 Mhz 时钟
always #10 clk = ~clk;

endmodule